module vcliargs

fn test_key() {
	
}
