module vcliargs

fn test_convert() {
	
}
