module vcliargs

fn test_parse() {

}
